-------------------------------------------------------------------------------------------------
-- Company   : CNES
-- Author    : John Doe (Developper Company JohnDoeCompany on behalf of ContractorBigcompany )
-- Copyright : Copyright (c) CNES.
-- Licensing : This VHDL entity can be licensed to be be used in the frame of CNES contracts.
--             Ask CNES for an end-user license agreement (EULA). 
-------------------------------------------------------------------------------------------------
-- Version         : V1
-- Version history : 
--    V1 : yyyy-mm-dd : Author name's John Doe (JohnDoeCompany): Creation
--    V2 : yyyy-mm-dd : Author name's John Toe (JohnToeCompany): 
--                         Modification description
--                         Modifications impacts
--                         Modifications reasons
-------------------------------------------------------------------------------------------------
-- File name          : header.vhd
-- File Creation date : yyyy-mm-dd
-- Project name       : VHDL Handbook CNES Edition 
-------------------------------------------------------------------------------------------------
-- Softwares             :  PC (OS version) - Editor (Version) - Synthetizer (Version) - P&R (Version)
-- Automatic VHDL coding :  YES/NO 
--                          Tool used + Version 
--                          Source file information
-------------------------------------------------------------------------------------------------
-- Description : Relevant information related to this entity 
--
-- Limitations : Hypothesis/constraints made on the external interfaces or configuration
--               that will impact this entity
--
-------------------------------------------------------------------------------------------------
-- Naming conventions: 
--
-- i_Port: Input entity port
-- o_Port: Output entity port
-- b_Port: Bidirectional entity port
-- g_My_Generic: Generic entity port
--
-- c_My_Constant: Constant definition 
-- t_My_Type: Custom type definition
--
-- My_Signal_n: Active low signal
-- v_My_Variable: Variable
-- sm_My_Signal: FSM signal
-- pkg_Param: Element Param coming from a package
--
-- My_Signal_re: Rising edge detection of My_Signal
-- My_Signal_fe: Falling edge detection of My_Signal
-- My_Signal_rX: X times registered My_Signal signal
--
-- P_Process_Name: Process
--
-------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity header is
    port  (

    );
end header;

architecture Behavioral of header is
begin
   -- Behavioral code of header
end Behavioral;